module demux ( 
	c,
	d,
	e,
	f,
	g,
	a,
	b,
	s,
	o
	) ;

input  c;
input  d;
input  e;
input  f;
input  g;
input  a;
input  b;
input [2:0] s;
inout  o;
